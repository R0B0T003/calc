module seven_seg(in, clr, seg1, seg2, seg3, seg4);
	input [7:0] in;
	input clr;
	output reg [6:0] seg1, seg2, seg3, seg4;
	wire [3:0] thos, huns, tens, unit;
	binary_to_bcd_converter bcd1(in, clr, unit, tens, huns, thos);
	
	
	always @(in, clr)
	begin
	case(thos)
		4'b0000 : seg4 = 7'b1000000; //0
		4'b0001 : seg4 = 7'b1111001; //1
		4'b0010 : seg4 = 7'b0100100; //2
		4'b0011 : seg4 = 7'b0110000; //3
		4'b0100 : seg4 = 7'b0011001; //4
		4'b0101 : seg4 = 7'b0010010; //5
		4'b0110 : seg4 = 7'b0000010; //6
		4'b0111 : seg4 = 7'b1111000; //7
		4'b1000 : seg4 = 7'b0000000; //8
		4'b1001 : seg4 = 7'b0010000; //9
		4'b1010 : seg4 = 7'b0001000; //A
		4'b1011 : seg4 = 7'b0000011; //b
		4'b1100 : seg4 = 7'b1000110; //C
		4'b1101 : seg4 = 7'b0100001; //D
		4'b1110 : seg4 = 7'b0000110; //E
		4'b1111 : seg4 = 7'b0001110; //F
		default : seg4 = 7'b1000000;
	endcase
	case(huns)
		4'b0000 : seg3 = 7'b1000000; //0
		4'b0001 : seg3 = 7'b1111001; //1
		4'b0010 : seg3 = 7'b0100100; //2
		4'b0011 : seg3 = 7'b0110000; //3
		4'b0100 : seg3 = 7'b0011001; //4
		4'b0101 : seg3 = 7'b0010010; //5
		4'b0110 : seg3 = 7'b0000010; //6
		4'b0111 : seg3 = 7'b1111000; //7
		4'b1000 : seg3 = 7'b0000000; //8
		4'b1001 : seg3 = 7'b0010000; //9
		4'b1010 : seg3 = 7'b0001000; //A
		4'b1011 : seg3 = 7'b0000011; //b
		4'b1100 : seg3 = 7'b1000110; //C
		4'b1101 : seg3 = 7'b0100001; //D
		4'b1110 : seg3 = 7'b0000110; //E
		4'b1111 : seg3 = 7'b0001110; //F
		default: seg3 = 7'b1000000;
	endcase		

		
	case(tens)
		4'b0000 : seg2 = 7'b1000000; //0
		4'b0001 : seg2 = 7'b1111001; //1
		4'b0010 : seg2 = 7'b0100100; //2
		4'b0011 : seg2 = 7'b0110000; //3
		4'b0100 : seg2 = 7'b0011001; //4
		4'b0101 : seg2 = 7'b0010010; //5
		4'b0110 : seg2 = 7'b0000010; //6
		4'b0111 : seg2 = 7'b1111000; //7
		4'b1000 : seg2 = 7'b0000000; //8
		4'b1001 : seg2 = 7'b0010000; //9
		4'b1010 : seg2 = 7'b0001000; //A
		4'b1011 : seg2 = 7'b0000011; //b
		4'b1100 : seg2 = 7'b1000110; //C
		4'b1101 : seg2 = 7'b0100001; //D
		4'b1110 : seg2 = 7'b0000110; //E
		4'b1111 : seg2 = 7'b0001110; //F
		default: seg2 = 7'b1000000;
	endcase		
	case(unit)
		4'b0000 : seg1 = 7'b1000000; //0
		4'b0001 : seg1 = 7'b1111001; //1
		4'b0010 : seg1 = 7'b0100100; //2
		4'b0011 : seg1 = 7'b0110000; //3
		4'b0100 : seg1 = 7'b0011001; //4
		4'b0101 : seg1 = 7'b0010010; //5
		4'b0110 : seg1 = 7'b0000010; //6
		4'b0111 : seg1 = 7'b1111000; //7
		4'b1000 : seg1 = 7'b0000000; //8
		4'b1001 : seg1 = 7'b0010000; //9
		4'b1010 : seg1 = 7'b0001000; //A
		4'b1011 : seg1 = 7'b0000011; //b
		4'b1100 : seg1 = 7'b1000110; //C
		4'b1101 : seg1 = 7'b0100001; //D
		4'b1110 : seg1 = 7'b0000110; //E
		4'b1111 : seg1 = 7'b0001110; //F
		default: seg1 = 7'b1000000;
	endcase
	
	end
		
		
endmodule 